package reg_seq_pkg;

import Registers_pkg::*;
import reg_model_pkg::*;
import shared_pkg::*;
import 
import uvm_pkg::*;
 `include "uvm_macros.svh"

 class reg_seq extends uvm_reg_sequence;
    function new();
        
    endfunction //new()
 endclass //reg_seq extends superClass

    
endpackage