`timescale 1ps/1ps
package Ram_config_pkg;
import shared_pkg::*;
import uvm_pkg::*;
`include "uvm_macros.svh"

// Configration class

endpackage