package shared_pkg;
    parameter ADDR_WIDTH = 32;
    parameter DATA_WIDTH = 32;
    parameter PSTRB_WIDTH = DATA_WIDTH/8;
    parameter ADDR_slave = 2'b00 ;
    parameter MY_PROT = 3'b000;
endpackage