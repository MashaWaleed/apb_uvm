package shared_pkg;
    parameter ADDR_WIDTH = 16;
    parameter DATA_WIDTH = 32;
    parameter PSTRB_WIDTH = DATA_WIDTH/8;
endpackage