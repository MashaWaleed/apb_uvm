package driver_pkg;
    import uvm_pkg::*;
    import shared_pkg::*;
    import config_pkg::*;

    `include "uvm_macros.svh"

    `include "apb_driver.sv"
    `include "uart_rx_driver.sv"
    `include "Ram_driver.sv"
endpackage