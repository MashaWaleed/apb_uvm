package sequenceItem_pkg;
    import uvm_pkg::*;
    import shared_pkg::*;
    import config_pkg::*;

    `include "uvm_macros.svh"

    `include "apb_sequence_item.sv"
    `include "uart_rx_sequence_item.sv"
    `include "Ram_sequenceItem.sv"

endpackage